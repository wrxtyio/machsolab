/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : logisimTopLevelShell                                         **
 **                                                                          **
 *****************************************************************************/

module logisimTopLevelShell( A_0,
                             B_0,
                             C_0 );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input A_0;
   input B_0;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output C_0;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire s_A;
   wire s_B;
   wire s_C;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** All signal adaptations are performed here                                  **
   *******************************************************************************/
   assign C_0 = s_C;
   assign s_A = A_0;
   assign s_B = B_0;

   /*******************************************************************************
   ** The toplevel component is connected here                                   **
   *******************************************************************************/
   test   CIRCUIT_0 (.A(s_A),
                     .B(s_B),
                     .C(s_C));
endmodule
